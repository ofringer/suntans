netcdf Estuary_IC {
dimensions:
	Nc = 4446 ;
	Np = 2348 ;
	Ne = 6793 ;
	Nk = 24 ;
	Nkw = 25 ;
	numsides = 3 ;
	two = 2 ;
	time = UNLIMITED ; // (1 currently)
variables:
	int suntans_mesh ;
		suntans_mesh:long_name = "Topology data of 2D unstructured mesh" ;
		suntans_mesh:edge_coordinates = "xe ye" ;
		suntans_mesh:face_edge_connectivity = "face" ;
		suntans_mesh:topology_dimension = "2" ;
		suntans_mesh:edge_face_connectivity = "grad" ;
		suntans_mesh:edge_node_connectivity = "edges" ;
		suntans_mesh:node_coordinates = "xp yp" ;
		suntans_mesh:cf_role = "mesh_topology" ;
		suntans_mesh:face_node_connectivity = "cells" ;
		suntans_mesh:face_coordinates = "xv yv" ;
	int cells(Nc, numsides) ;
		cells:long_name = "Maps every face to its corner nodes" ;
		cells:cf_role = "face_node_connectivity" ;
	int edges(Ne, two) ;
		edges:long_name = "Maps every edge to the two nodes it connects" ;
		edges:cf_role = "edge_node_connectivity" ;
	int neigh(Nc, numsides) ;
		neigh:long_name = "Maps every face to its neighbouring faces" ;
		neigh:cf_role = "face_face_connectivity" ;
	int grad(Ne, two) ;
		grad:long_name = "Maps every edge to the two faces it connects" ;
		grad:cf_role = "edge_face_connectivity" ;
	double xp(Np) ;
		xp:long_name = "Easting of 2D mesh node" ;
		xp:standard_name = "Easting" ;
	double yp(Np) ;
		yp:long_name = "Northing of 2D mesh nodes" ;
		yp:standard_name = "Northing" ;
	double xv(Nc) ;
		xv:long_name = "Easting of 2D mesh face" ;
		xv:standard_name = "Easting" ;
	double yv(Nc) ;
		yv:long_name = "Easting of 2D mesh face" ;
		yv:standard_name = "Easting" ;
	double dv(Nc) ;
		dv:positive = "down" ;
		dv:coordinates = "xv yv" ;
		dv:long_name = "seafloor depth" ;
		dv:standard_name = "sea_floor_depth_below_geoid" ;
		dv:mesh = "suntans_mesh" ;
		dv:location = "face" ;
		dv:units = "m" ;
	double dz(Nk) ;
		dz:units = "m" ;
		dz:long_name = "z layer spacing" ;
	double z_r(Nk) ;
		z_r:units = "m" ;
		z_r:long_name = "depth at layer mid points" ;
		z_r:standard_name = "ocean_z_coordinate" ;
		z_r:positive = "up" ;
	int Nk(Nc) ;
		Nk:long_name = "Number of layers at face" ;
	double time(time) ;
		time:_FillValue = 999999. ;
		time:units = "seconds since 1990-01-01 00:00:00" ;
		time:long_name = "time" ;
	double eta(time, Nc) ;
		eta:_FillValue = 999999. ;
		eta:units = "metres" ;
		eta:long_name = "Sea surface elevation" ;
	double uc(time, Nk, Nc) ;
		uc:_FillValue = 999999. ;
		uc:units = "metre second-1" ;
		uc:long_name = "Eastward water velocity component" ;
	double vc(time, Nk, Nc) ;
		vc:_FillValue = 999999. ;
		vc:units = "metre second-1" ;
		vc:long_name = "Northward water velocity component" ;
	double S(time, Nk, Nc) ;
		S:_FillValue = 999999. ;
		S:units = "ppt" ;
		S:long_name = "Salinity" ;
	double T(time, Nk, Nc) ;
		T:_FillValue = 999999. ;
		T:units = "degrees C" ;
		T:long_name = "Water temperature" ;

// global attributes:
		:Description = "SUNTANS History file" ;
		:Author = "" ;
		:Created = "2013-04-09T09:35:25.094231" ;
}
