netcdf Estuary_BC {
dimensions:
	Nt = UNLIMITED ; // (1465 currently)
	Nk = 24 ;
	Ntype2 = 7 ;
	Ntype3 = 77 ;
	Nseg = 1 ;
variables:
	double xv(Ntype3) ;
		xv:long_name = "Easting of type-3 boundary points" ;
		xv:units = "metres" ;
	double yv(Ntype3) ;
		yv:long_name = "Northing of type-3 boundary points" ;
		yv:units = "metres" ;
	int cellp(Ntype3) ;
		cellp:long_name = "Index of suntans grid cell corresponding to type-3 boundary" ;
		cellp:units = "" ;
	double xe(Ntype2) ;
		xe:long_name = "Easting of type-2 boundary points" ;
		xe:units = "metres" ;
	double ye(Ntype2) ;
		ye:long_name = "Northing of type-2 boundary points" ;
		ye:units = "metres" ;
	int edgep(Ntype2) ;
		edgep:long_name = "Index of suntans grid edge corresponding to type-2 boundary" ;
		edgep:units = "" ;
	int segedgep(Ntype2) ;
		segedgep:long_name = "Pointer to boundary segment flag for each type-2 edge" ;
		segedgep:units = "" ;
	int segp(Nseg) ;
		segp:long_name = "Boundary segment flag" ;
		segp:units = "" ;
	double z(Nk) ;
		z:long_name = "Vertical grid mid-layer depth" ;
		z:units = "metres" ;
	double time(Nt) ;
		time:long_name = "Boundary time" ;
		time:units = "seconds since 1990-01-01 00:00:00" ;
	double boundary_u(Nt, Nk, Ntype2) ;
		boundary_u:long_name = "Eastward velocity at type-2 boundary point" ;
		boundary_u:units = "metre second-1" ;
	double boundary_v(Nt, Nk, Ntype2) ;
		boundary_v:long_name = "Northward velocity at type-2 boundary point" ;
		boundary_v:units = "metre second-1" ;
	double boundary_w(Nt, Nk, Ntype2) ;
		boundary_w:long_name = "Vertical velocity at type-2 boundary point" ;
		boundary_w:units = "metre second-1" ;
	double boundary_T(Nt, Nk, Ntype2) ;
		boundary_T:long_name = "Water temperature at type-2 boundary point" ;
		boundary_T:units = "degrees C" ;
	double boundary_S(Nt, Nk, Ntype2) ;
		boundary_S:long_name = "Salinity at type-2 boundary point" ;
		boundary_S:units = "psu" ;
	double boundary_Q(Nt, Nseg) ;
		boundary_Q:long_name = "Volume flux  at boundary segment" ;
		boundary_Q:units = "metre^3 second-1" ;
	double uc(Nt, Nk, Ntype3) ;
		uc:long_name = "Eastward velocity at type-3 boundary point" ;
		uc:units = "metre second-1" ;
	double vc(Nt, Nk, Ntype3) ;
		vc:long_name = "Northward velocity at type-3 boundary point" ;
		vc:units = "metre second-1" ;
	double wc(Nt, Nk, Ntype3) ;
		wc:long_name = "Vertical velocity at type-3 boundary point" ;
		wc:units = "metre second-1" ;
	double T(Nt, Nk, Ntype3) ;
		T:long_name = "Water temperature at type-3 boundary point" ;
		T:units = "degrees C" ;
	double S(Nt, Nk, Ntype3) ;
		S:long_name = "Salinity at type-3 boundary point" ;
		S:units = "psu" ;
	double h(Nt, Ntype3) ;
		h:long_name = "Water surface elevation at type-3 boundary point" ;
		h:units = "metres" ;
}
