netcdf Estuary_MetForcing {
dimensions:
	nt = UNLIMITED ; // (1465 currently)
	NUwind = 1 ;
	NVwind = 1 ;
	NTair = 1 ;
	NPair = 1 ;
	NRH = 1 ;
	Nrain = 1 ;
	Ncloud = 1 ;
variables:
	double Time(nt) ;
		Time:long_name = "time" ;
		Time:units = "seconds since 1990-01-01 00:00:00" ;
	double x_Uwind(NUwind) ;
		x_Uwind:long_name = "Longitude at Uwind" ;
		x_Uwind:units = "degrees_north" ;
	double y_Uwind(NUwind) ;
		y_Uwind:long_name = "Latitude at Uwind" ;
		y_Uwind:units = "degrees_east" ;
	double z_Uwind(NUwind) ;
		z_Uwind:long_name = "Elevation at Uwind" ;
		z_Uwind:units = "m" ;
	double x_Vwind(NVwind) ;
		x_Vwind:long_name = "Longitude at Vwind" ;
		x_Vwind:units = "degrees_north" ;
	double y_Vwind(NVwind) ;
		y_Vwind:long_name = "Latitude at Vwind" ;
		y_Vwind:units = "degrees_east" ;
	double z_Vwind(NVwind) ;
		z_Vwind:long_name = "Elevation at Vwind" ;
		z_Vwind:units = "m" ;
	double x_Tair(NTair) ;
		x_Tair:long_name = "Longitude at Tair" ;
		x_Tair:units = "degrees_north" ;
	double y_Tair(NTair) ;
		y_Tair:long_name = "Latitude at Tair" ;
		y_Tair:units = "degrees_east" ;
	double z_Tair(NTair) ;
		z_Tair:long_name = "Elevation at Tair" ;
		z_Tair:units = "m" ;
	double x_Pair(NPair) ;
		x_Pair:long_name = "Longitude at Pair" ;
		x_Pair:units = "degrees_north" ;
	double y_Pair(NPair) ;
		y_Pair:long_name = "Latitude at Pair" ;
		y_Pair:units = "degrees_east" ;
	double z_Pair(NPair) ;
		z_Pair:long_name = "Elevation at Pair" ;
		z_Pair:units = "m" ;
	double x_RH(NRH) ;
		x_RH:long_name = "Longitude at RH" ;
		x_RH:units = "degrees_north" ;
	double y_RH(NRH) ;
		y_RH:long_name = "Latitude at RH" ;
		y_RH:units = "degrees_east" ;
	double z_RH(NRH) ;
		z_RH:long_name = "Elevation at RH" ;
		z_RH:units = "m" ;
	double x_rain(Nrain) ;
		x_rain:long_name = "Longitude at rain" ;
		x_rain:units = "degrees_north" ;
	double y_rain(Nrain) ;
		y_rain:long_name = "Latitude at rain" ;
		y_rain:units = "degrees_east" ;
	double z_rain(Nrain) ;
		z_rain:long_name = "Elevation at rain" ;
		z_rain:units = "m" ;
	double x_cloud(Ncloud) ;
		x_cloud:long_name = "Longitude at cloud" ;
		x_cloud:units = "degrees_north" ;
	double y_cloud(Ncloud) ;
		y_cloud:long_name = "Latitude at cloud" ;
		y_cloud:units = "degrees_east" ;
	double z_cloud(Ncloud) ;
		z_cloud:long_name = "Cloud cover fraction" ;
		z_cloud:units = "Fraction (0-1)" ;
	double Uwind(nt, NUwind) ;
		Uwind:coordinates = "x_Uwind,y_Uwind" ;
	double Vwind(nt, NVwind) ;
		Vwind:coordinates = "x_Vwind,y_Vwind" ;
	double Tair(nt, NTair) ;
		Tair:coordinates = "x_Tair,y_Tair" ;
	double Pair(nt, NPair) ;
		Pair:coordinates = "x_Pair,y_Pair" ;
	double RH(nt, NRH) ;
		RH:coordinates = "x_RH,y_RH" ;
	double rain(nt, Nrain) ;
		rain:coordinates = "x_rain,y_rain" ;
	double cloud(nt, Ncloud) ;
		cloud:coordinates = "x_cloud,y_cloud" ;
}
